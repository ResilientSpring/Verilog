`timescale 50ps/1ps

module light2(x1, x2, f);

input x1, x2;
output f;



endmodule