module BlinkLEDs1 (
    Clock, Reset, OUT_High, OUT_low
);

input Clock, Reset;
output OUT_High, OUT_low;
    
endmodule