module TopLevel (
    // names for pins  
    // each name represents a pin or a vector of pins
    SW,
    LEDR
);

input [0:9] SW;
output 
    
endmodule