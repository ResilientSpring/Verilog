module TopLevel (
    SW, LEDR, HEX0, HEX1, HEX2, HEX3
);

input [9:0] SW;
output [9:0] LEDR;
output [7:0] HEX0, HEX1, HEX2, HEX3;


    
endmodule