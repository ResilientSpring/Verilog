// Verilog arithmetic operator

module arithmetic_operation (a, b, y1, y2, y3, y4, y5);

input [0:3] a, b;
output [0:4] y1;
output [0:5] y3;
output [0:3] y2, y4, y5;



endmodule