module Logic_optimization (
    a, b, c, d, m, n
);

input a, b, c, d;
output m, n;

and ac(a, c);

    
endmodule