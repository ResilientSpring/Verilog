module TopLevel (
    input [1:0] SW,
    output [1:0] LEDR
);



always @(*) begin


end

    
endmodule