module TopLevel (
    input [0:5] SW,
    output [0:5] LEDR,
    output HEX0, HEX1, HEX2, HEX3, HEX4, HEX5
);


    
endmodule