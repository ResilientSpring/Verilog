module first_system (
    out1, out2, in1, in2
);

// Port definitions
input in1, in2;
output out1, out2;

// Description of the digital system
// Dataflow modeling

wire and_out, or_out;

    
endmodule