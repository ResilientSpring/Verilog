module TopLevel (
    input [9:0] SW, 
    output [9:0] LEDR
);
    
endmodule