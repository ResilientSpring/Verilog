module TopLevel (
    SW, LEDR
);

input [9:0] SW;
output [9:0] LEDR;
    
endmodule