module  (
    switches,
    HEXo
);

input [0:6] switches;
output [0:6] HEXo;

    
endmodule