module TopLevel (
    // names for pins  
    // (Each name can represent a single pin or a vector - group of pins)
    SW,
    LEDR
);

input [0:9] SW;
output 
    
endmodule