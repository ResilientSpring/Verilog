module TopLevel (
    SW,
    LEDR,
    HEX0,, HEX1, HEX2, HEX3, HEX4, HEX5
);
    
    


endmodule